module decrypt#(parameter nk=4,parameter nr=10)(input [0:127]in ,output [0:127]out,input [0:128*(nr+1)-1] key_d);  // nb*(nr+1) words where nb always = 4 and 1 word = 4 bytes = 32 bit so 32*4=128

endmodule